module Mineswepper (
input [3:0] kb_row, kb_col, // keyboard
input CLK,
output A,B,C,D,E,F,G // 7 seg
);
















endmodule